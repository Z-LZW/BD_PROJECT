`ifndef SYSTEM_INTERFACE_GUARD
`define SYSTEM_INTERFACE_GUARD

interface system_interface(output bit clk, rst_n);
endinterface

`endif