`include "base_test.sv"
`include "register_sanity_test.sv"
`include "basic_master_read_test.sv"
`include "basic_master_write_test.sv"
`include "fifo_full_test.sv"
`include "basic_slave_rx_test.sv"
`include "basic_slave_tx_test.sv"