`ifndef CONF_MASTER_WRITE_GUARD
`define CONF_MASTER_WRITE_GUARD

class configure_master_write extends virtual_sequence_base;
  
  uvm_status_e status;
  uvm_reg_data_t data;

  //address register
  rand bit [7-1:0] target_addr;

  //control register
  rand bit [8-1:0] tx_lim    ;

  //irq mask register
  rand bit         rx_fifo_empty_mask;
  rand bit         tx_fifo_full_mask;
  rand bit         rx_fail_mask;
  rand bit         tx_fail_mask;
  rand bit         rx_done_mask;
  rand bit         tx_done_mask;

  rand bit         read;

  //divider
  rand bit [16-1:0] divider;

  `uvm_object_utils(configure_master_write)   

  function new(string name = "configure_master_write");
    super.new(name);
  endfunction:new 

  function randomize();
    assert (std::randomize(target_addr)) else $fatal("randomization failed in master write configuration sequence");

    assert (std::randomize(tx_lim)) else $fatal("randomization failed in master write configuration sequence");

    assert (std::randomize(rx_fifo_empty_mask)) else $fatal("randomization failed in master write configuration sequence");
    assert (std::randomize(tx_fifo_full_mask)) else $fatal("randomization failed in master write configuration sequence");
    assert (std::randomize(rx_fail_mask)) else $fatal("randomization failed in master write configuration sequence");
    assert (std::randomize(tx_fail_mask)) else $fatal("randomization failed in master write configuration sequence");
    assert (std::randomize(rx_done_mask)) else $fatal("randomization failed in master write configuration sequence");
    assert (std::randomize(tx_done_mask)) else $fatal("randomization failed in master write configuration sequence");

    assert (std::randomize(read)) else $fatal("randomization failed in master write configuration sequence");

    assert (std::randomize(divider)) else $fatal("randomization failed in master write configuration sequence");
  endfunction

  virtual task body();
    p_sequencer.p_reg_model.divider.write(status,divider);              //set divider
    p_sequencer.p_reg_model.ctrl.write(status,{tx_lim,5'b0,'h7});       //set transfer limit | enable device | enable ack | mode
    p_sequencer.p_reg_model.cmd.write(status,'h1c);                     //clear the interrupt and fifos
    p_sequencer.p_reg_model.addr.write(status,{target_addr,8'b0});      //write the target address

    repeat(tx_lim) begin
      p_sequencer.p_reg_model.tx_fifo_data.write(status,data);          //write the data in the tx fifo
    end

    p_sequencer.p_reg_model.irq_mask.write(status,{rx_fifo_empty_mask,
                                                   rx_fifo_empty_mask,
                                                   rx_fail_mask,
                                                   tx_fail_mask,
                                                   rx_done_mask,
                                                   tx_done_mask});      //masking the coresponding interrupts

    p_sequencer.p_reg_model.cmd.write(status,{read,1'b1});              //initiate write
      
  endtask
endclass

`endif