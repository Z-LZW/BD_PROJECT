`ifndef APB_PACKAGE_GUARD
`define APB_PACKAGE_GUARD

package apb_package
  
  import uvm_pkg::*;

  `include "apb_if.sv"
  `include "apb_types.sv"
  `include "apb_trans.sv"
  `include "apb_diver.sv"
  `include "apb_monitor.sv"
  `include "apb_base_sequence.sv"
  `include "apb_sequencer.sv"
  `include "apb_coverage.sv"
  `include "apb_agent.sv"

endpackage

`endif