`include "base_test.sv"
`include "apb_selfcheck.sv"
`include "i2c_selfcheck.sv"