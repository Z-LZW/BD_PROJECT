`ifndef APB_PACKAGE_GUARD
`define APB_PACKAGE_GUARD

package apb_package;
  
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "apb_types.sv"
  `include "apb_trans.sv"
  `include "apb_driver.sv"
  `include "apb_monitor.sv"
  //`include "apb_base_sequence.sv"
  `include "apb_sequencer.sv"
  `include "apb_coverage.sv"
  `include "apb_agent.sv"

endpackage

`endif