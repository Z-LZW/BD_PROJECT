`include "configure_master_read.sv"
`include "configure_master_write.sv"
`include "configure_slave.sv"
`include "i2c_master_read_seq.sv"
`include "i2c_master_write_seq.sv"
`include "i2c_slave_seq.sv"
`include "poll_status.sv"
`include "read_every_register.sv"
`include "read_irq.sv"
`include "read_rx_fifo.sv"
`include "system_reset_sequence.sv"
`include "write_every_register.sv"
