`ifndef SYSTEM_PACKAGE_GUARD
`define SYSTEM_PACKAGE_GUARD

package system_package;

  `include "system_if.sv"
  `include "system_trans.sv"

endpackage

`endif 